-- Implement the architecture for the game here (Exercise II)
