
library ieee;
use ieee.std_logic_1164.all;

package gfx_init_pkg is
	type gfx_init_cmds_t is array(natural range<>) of std_logic_vector;
	
	constant GFX_INIT_CMDS : gfx_init_cmds_t(0 to 1725) := (
	x"9000",
	x"0000",
	x"0000",
	x"0140",
	x"00f0",
	x"9001",
	x"2c00",
	x"0001",
	x"0140",
	x"00f0",
	x"9002",
	x"5800",
	x"0002",
	x"0158",
	x"0008",
	x"7001",
	x"0560",
	x"5800",
	x"0002",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"00ff",
	x"ff00",
	x"ffff",
	x"0000",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"0000",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"0000",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"9003",
	x"62c0",
	x"0002",
	x"0050",
	x"0008",
	x"7001",
	x"0140",
	x"62c0",
	x"0002",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ff00",
	x"00ff",
	x"ff00",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"00ff",
	x"ff00",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ff00",
	x"0000",
	x"0000",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"0000",
	x"00ff",
	x"ff00",
	x"0000",
	x"00ff",
	x"ff00",
	x"00ff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ff00",
	x"00ff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"ffff",
	x"0000",
	x"00ff",
	x"ff00",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"00ff",
	x"ff00",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ff00",
	x"00ff",
	x"ff00",
	x"00ff",
	x"0000",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"0000",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ff00",
	x"00ff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"ffff",
	x"ffff",
	x"00ff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ffff",
	x"ff00",
	x"ffff",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"0000",
	x"ff00",
	x"ffff",
	x"8000",
	x"84ff"
	);
end package;

