-- put your implementation the dualshock_ctrl here (Exercise II)
